library ieee;
use ieee.std_logic_1164.all;

entity rom is
	generic( n : integer := 64 ); 		 -- tama�o de palabra
	port(
		m1,m2,b1,b2,a,x0: out	std_logic_vector(n-1 downto 0)
	);	
end rom;					 

architecture arch of rom is
begin	  	
 m1 <= "0000000001100110011001100110011001100110011001100110011001101000";	 --      0.800 
 m2 <= "0000001010000000000000000000000000000000000000000000000000000000";	 --      5.000 
 b1 <= "0000001000000000000000000000000000000000000000000000000000000000";	 --      4.000 
 b2 <= "0000110010000000000000000000000000000000000000000000000000000000";	 --     25.000 
  a <= "0000001010000000000000000000000000000000000000000000000000000000";	 --      5.000 
 x0 <= "0000000000001100110011001100110011001100110011001100110011001101";	 --      0.100
	 
	 
end arch;
